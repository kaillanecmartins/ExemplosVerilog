// Aula 01 - Exemplos
module porta_not(
	input a,
  	output y
);
  
  assign y = ~a;
endmodule