// Aula 01 - Exemplos
module porta_and(
	input a,
  	input b,
  	output y
);
  
  assign y = a & b;
endmodule